----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Izel Molina & Brandan Jimenez
-- 
-- Create Date: 26.02.2021 19:51:41
-- Design Name: Alarm
-- Module Name: Alarm - Behavioral
-- Project Name: Practica 5
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Alarm is
        Port(clk_input: in bit;
            PM: out bit);
            --input: in bit := '1';
            --hrs_dec, AM, PM: out bit;
            --hrs_uni, min_uni, seg_uni: out bit_vector(3 downto 0);
            --min_dec, seg_dec: out bit_vector(2 downto 0));
end Alarm;

architecture Behavioral of Alarm is
    
    component FFJK
        Port(J, K, resetN, setN, clk: in bit;
            Q, Qnot: out bit);
    end component;
    
    component CounterHrsMOD12
        Port(clk: in bit;
            input: in bit:= '1';
            hrs_uni: out bit_vector(3 downto 0);
            hrs_dec: out bit);
    end component;
    
    component CounterMinMOD60
        Port(clk, input: in bit;
             min_uni: out bit_vector(3 downto 0);
             min_dec: out bit_vector(2 downto 0));
    end component;
    
    component CounterSecMOD60
        Port(clk, input: in bit;
            seg_uni: out bit_vector(3 downto 0);
            seg_dec: out bit_vector(2 downto 0));
    end component;
    
    component sSegDisplay is
        Port(ck : in  bit;                          -- 100MHz system clock
                number : in  bit_vector (63 downto 0); -- eight digit number to be displayed
                seg : out  bit_vector (7 downto 0);    -- display cathodes
                an : out  bit_vector (7 downto 0));    -- display anodes (active-low, due to transistor complementing)
    end component;

signal input: bit := '1';
signal clk_divisor: integer := 0;
signal startHrsCounter, AM_PM, AM, internal_hrs_dec, clk_in: bit;
signal internal_min_dec, internal_sec_dec: bit_vector(2 downto 0);
signal internal_hrs_uni, internal_min_uni, internal_sec_uni: bit_vector(3 downto 0);
signal d7s: bit_vector(63 downto 0) := "1111111111111111111111111111111100000000000000000000000000000000";  

begin
    process(clk_in, clk_input)
    begin
    --A�adir el divisor de frecuencia 1x10^8
        if clk_input'event and clk_input = '1' then
           divisor: if clk_divisor <= 50000000 then
                --wait until clk_input'event and clk_input = '1';
                clk_divisor <= clk_divisor + 1;
                if clk_divisor = 100000000 then
                    clk_in <= '1';
                    clk_divisor <= 0;
                else
                    clk_in <= '0';
                end if;    
            end if;
          end if;
         
        if CLK_IN'event and clk_in = '1' then
            startHrsCounter <=  internal_min_dec(2) and internal_min_dec(0) and internal_min_uni(3) and internal_min_uni(0) and 
                                internal_sec_dec(2) and internal_sec_dec(0) and internal_sec_uni(3) and internal_sec_uni(0); 
                                    
            AM_PM           <=  internal_hrs_dec and internal_hrs_uni(0) and internal_min_dec(2) and internal_min_dec(0) and internal_min_uni(3) 
                                and internal_min_uni(0) and internal_sec_dec(2) and internal_sec_dec(0) and internal_sec_uni(3) and internal_sec_uni(0); 
        end if;
    
        case (internal_min_uni) is
                        when "0000" => d7s(15 downto 8) <= "11000000";
                        when "0001" => d7s(15 downto 8) <= "11111001";
                        when "0010" => d7s(15 downto 8) <= "10100100";
                        when "0011" => d7s(15 downto 8) <= "10110000";
                        when "0100" => d7s(15 downto 8) <= "10011001";
                        when "0101" => d7s(15 downto 8) <= "10010010";
                        when "0110" => d7s(15 downto 8) <= "10000010";
                        when "0111" => d7s(15 downto 8) <= "11111000";
                        when "1000" => d7s(15 downto 8) <= "10000000";
                        when "1001" => d7s(15 downto 8) <= "10010000";
                        when others => d7s(15 downto 8) <= "11111111";
                        end case;
         
        case (internal_hrs_uni) is
                        when "0000" => d7s(15 downto 8) <= "11000000";
                        when "0001" => d7s(15 downto 8) <= "11111001";
                        when "0010" => d7s(15 downto 8) <= "10100100";
                        when "0011" => d7s(15 downto 8) <= "10110000";
                        when "0100" => d7s(15 downto 8) <= "10011001";
                        when "0101" => d7s(15 downto 8) <= "10010010";
                        when "0110" => d7s(15 downto 8) <= "10000010";
                        when "0111" => d7s(15 downto 8) <= "11111000";
                        when "1000" => d7s(15 downto 8) <= "10000000";
                        when "1001" => d7s(15 downto 8) <= "10010000";
                        when others => d7s(15 downto 8) <= "11111111";
                        end case;
            
        case (internal_min_dec) is
                        when "000" => d7s(15 downto 8) <= "11000000";
                        when "001" => d7s(15 downto 8) <= "11111001";
                        when "010" => d7s(15 downto 8) <= "10100100";
                        when "011" => d7s(15 downto 8) <= "10110000";
                        when "100" => d7s(15 downto 8) <= "10011001";
                        when "101" => d7s(15 downto 8) <= "10010010";
                        --when "0110" => d7s(15 downto 8) <= "10000010";
                        --when "0111" => d7s(15 downto 8) <= "11111000";
                        --when "1000" => d7s(15 downto 8) <= "10000000";
                        --when "1001" => d7s(15 downto 8) <= "10010000";
                        when others => d7s(15 downto 8) <= "11111111";
                        end case;
        
        case (internal_hrs_dec) is
                        when '0' => d7s(15 downto 8) <= "11000000";
                        when '1' => d7s(15 downto 8) <= "11111001";
                        --when "010" => d7s(15 downto 8) <= "10100100";
                        --when "011" => d7s(15 downto 8) <= "10110000";
                        --when "100" => d7s(15 downto 8) <= "10011001";
                        --when "101" => d7s(15 downto 8) <= "10010010";
                        --when "0110" => d7s(15 downto 8) <= "10000010";
                        --when "0111" => d7s(15 downto 8) <= "11111000";
                        --when "1000" => d7s(15 downto 8) <= "10000000";
                        --when "1001" => d7s(15 downto 8) <= "10010000";
                        when others => d7s(15 downto 8) <= "11111111";
                        end case;
    end process; 
       
    --seg_uni <= internal_sec_uni;
    --seg_dec <= internal_sec_dec;
    --min_uni <= internal_min_uni;
    --min_dec <= internal_min_dec;
    --hrs_uni <= internal_hrs_uni;
    --hrs_dec <= internal_hrs_dec;
    
    CSM60:  CounterSecMOD60 port map (clk_in, input, internal_sec_uni, internal_sec_dec);
    CMM60:  CounterMinMOD60 port map (clk_in, input, internal_min_uni, internal_min_dec);
    CHM12:  CounterHrsMOD12 port map (startHrsCounter, input, internal_hrs_uni, internal_hrs_dec);
    AMPM:   FFJK port map (input, input, '1', '1', AM_PM, PM, AM);
end Behavioral;
